// lookup table
// deep 
// 9 bits wide; as deep as you wish
module InstrRom #(parameter D=9)(
  input       [D-1:0] prog_ctr,    // prog_ctr	  address pointer
  output logic[ 8:0] mach_code);

  logic[8:0] core[2**D];
  initial							    // load the program
  $readmemb("machine_code.txt",core);
  

  always_comb  begin
    mach_code = core[prog_ctr];
  end

endmodule


/*
sample mach_code.txt:

001111110		 // ADD r0 r1 r0
001100110
001111010
111011110
101111110
001101110
001000010
111011110
*/